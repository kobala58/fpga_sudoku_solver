module tb;
  test dut();
  initial begin
    #1;
    $finish;
  end
endmodule
